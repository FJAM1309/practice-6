module receiver (
);

endmodule 